module FA(input a, input b, input cin, output sum, output cout);
	wire w1, w2, w3;
	xor(w1, a, b);
	and(w2, a, b);
	xor(sum, w1, cin);
	and(w3, w1, cin);
	or(cout, w2, w3);
endmodule